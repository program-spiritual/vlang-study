module main

my_int := 1

my_closure := fn [my_int] () {
	println(my_int)
}

my_closure()

func :=fn[i]() int{
  return i
}

 println(func(1)==1)
 i=123
 println(func()==1)
