module main

import mymoudle2

fn main() {
	mymoudle2.say_hi()
	mymoudle2.say_hi_and_bye()
}
