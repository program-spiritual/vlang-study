module main

import sample

fn main() {
	println('Hello, World!')
	info := sample.new_information('sample information')!
	println(info)
}
